module calendar

pub struct Calendar {}
