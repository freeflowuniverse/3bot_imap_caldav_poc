module files

pub struct Files {}
